LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;


ENTITY test_comp IS

END ENTITY;

ARCHITECTURE test OF test_comp IS

COMPONENT n_bit_comparator IS
    GENERIC (length : INTEGER := 4);
    PORT (  a,b : IN STD_LOGIC_VECTOR(length-1 DOWNTO 0);
    led_upper,led_less,led_correct : OUT STD_LOGIC := 'Z');
END COMPONENT;

SIGNAL x,y                  : STD_LOGIC_vector(3 DOWNTO 0); 
SIGNAL UPPER,LESS,EQUAL     : STD_LOGIC;


BEGIN
    Stage : n_bit_comparator PORT MAP (x,y,UPPER,LESS,EQUAL);
    x  <= X"1",X"5" AFTER 200 NS,X"2" AFTER 400 NS,X"A" AFTER 600 NS; 
    y  <= X"2",X"4" AFTER 200 NS,X"2" AFTER 400 NS,X"F" AFTER 600 NS; 

END ARCHITECTURE;