LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Main IS

END ENTITY;

-----------------------------------------------------
-----------------------------------------------------
-----------------------------------------------------

ARCHITECTURE Main_ARCH OF Main IS
------------------------------------DECLARATION BEGIN


--------------------------------------END DECLARATION
BEGIN

END ARCHITECTURE;