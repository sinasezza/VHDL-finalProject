LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;


ENTITY seven_segment_tb IS

END ENTITY;


ARCHITECTURE test OF seven_segment_tb IS

COMPONENT seven_segment IS
    PORT(   threeBITinput  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
            eightBIToutput : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT;
SIGNAL  num     : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL  result  : STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
    mySTAGE : seven_segment PORT MAP(num,result);
    num <= "000" , "001" AFTER 100 NS , "010" AFTER 200 NS , "110" AFTER 400 ns;
END ARCHITECTURE;